module mux4ne1(
	input Hyrja0,
	input Hyrja1,
	input Hyrja2,
	input Hyrja3,
	input [1:0] S,
	output Dalja
	);
	assign Dalja =s[1] ? (S[0] ?Hyrja3 :Hyrja2) : (S[0] ? Hyrja1 :Hyrja0);
	
	endmodule 
	
	
